`ifndef __GLOBALS__
`define __GLOBALS__

// UVM Globals
localparam string IQ_IN_NAME = "1.0_read_IQ_output.txt";
localparam string LEFT_OUT_NAME = "uvm_leftout.txt";
localparam string RIGHT_OUT_NAME = "uvm_rightout.txt";
localparam string RIGHT_CMP_NAME = "2.8_out_right.txt";
localparam string LEFT_CMP_NAME = "1.8_out_left.txt";
localparam int CLOCK_PERIOD = 10;

`endif
